module main;
  initial
    begin
      $display("Alix(SenPai) - With love from Kavar Shiraz, IRAN");
      $finish;
    end
endmodule
